--------------------------------------------------------------------------------
--! @file
--! @brief XOROSHIRO128+ uniform random number generator
--! @author David Winter (adaption of the public domain XOROSHIRO128+)
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity xoroshiro128plus is
  generic (
    seed_1 : unsigned(63 downto 0);            --! first seed
    seed_0 : unsigned(63 downto 0)             --! second seed
    );
  port (
    clk    : in  std_logic;                    --! clock
    rstn   : in  std_logic;                    --! negative reset
    enable : in  std_logic;                    --! enable
    dout   : out std_logic_vector(63 downto 0) --! 64 bit uniform output
    );

end entity;

architecture beh of xoroshiro128plus is
  signal s_0 : std_logic_vector(63 downto 0);
  signal s_1 : std_logic_vector(63 downto 0);
begin

  dout <= std_logic_vector(unsigned(s_0) + unsigned(s_1));

  ctrl : process (clk, rstn)
    variable s_1n : std_logic_vector(63 downto 0);
  begin
    if rstn = '0' then
      s_0 <= std_logic_vector(seed_0);
      s_1 <= std_logic_vector(seed_1);
    elsif rising_edge(clk) and enable = '1' then
      s_1n := s_1 xor s_0;
      s_0  <= std_logic_vector((unsigned(s_0) rol 24) xor unsigned(s_1n) xor (unsigned(s_1n) sll 16));
      s_1  <= std_logic_vector(unsigned(s_1n) rol 37);
    end if;
  end process ctrl;

end architecture beh;


library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package xoro_seeds is
    type xoro_seed_t is array(1 downto 0) of unsigned(63 downto 0);
    type xoro_seeds_t is array(0 to 255) of xoro_seed_t;
    constant xoro_seeds : xoro_seeds_t := ((X"1976c51ab89a5886", X"86114fc94d6c4ad5"),
        (X"e0296ce69151a79f", X"99ee2d06176445b6"),
        (X"423716dc01d203b8", X"ead8937999d6599e"),
        (X"b23bc3269b334182", X"615f334a56ed3d96"),
        (X"f2ef604b534875ef", X"a5636f712dea8e2a"),
        (X"c3691e1ed3eba4ba", X"cfe05cb256d80bea"),
        (X"bedce2c93c1ea677", X"fa88764aca9d7688"),
        (X"0affa462a42fde70", X"4a64bd37250b762a"),
        (X"b8641e5cff3daf31", X"7a5501e6eca23cef"),
        (X"21d0edb5bbdd0eb2", X"61157fdec1979a79"),
        (X"c57fcc63470849a5", X"ba60076ce9ae3680"),
        (X"92e779b6933cd4f9", X"a24146171780a69c"),
        (X"a83cbdb0b9f3c874", X"08c56f09c31e7eff"),
        (X"192e0dd29ad9122e", X"c86d18a5e228a7e5"),
        (X"12f62825150f4826", X"44102a9b41b640b1"),
        (X"f59d7bd4f0f25b98", X"fbd060f2c2c89078"),
        (X"72eef6ecf3ee3408", X"17bf02e175df96f6"),
        (X"82607ac8844a0d0c", X"1de6e8268186f757"),
        (X"3276d8944cf53269", X"0c08d820c93bbafc"),
        (X"c72a56ea28195eb6", X"2390edd23f68a681"),
        (X"615eb1af63fcc0a1", X"553b6916a3621095"),
        (X"ff7c7809d00d28ca", X"1bee4a66f18702ee"),
        (X"aef96cc7087436d8", X"8fdddc3c43d88834"),
        (X"32e7ff4581fd9907", X"ca468296c56b0b55"),
        (X"a0c21eb30f847571", X"c44480d6df22eb96"),
        (X"ab76330cd68023b5", X"4641f041c2386626"),
        (X"29bdbf695f135db9", X"23ee7d29af119192"),
        (X"a5591829862caa8c", X"402e77bd8ebd6340"),
        (X"1ebc9a09f306eaa3", X"fd107eb4676626f0"),
        (X"fab275b8cceebce5", X"b57e6f5f6963fbbb"),
        (X"af2729c08939be92", X"9c47a631b3b820f9"),
        (X"acb38a17203b0b9e", X"06f15bea57b196ad"),
        (X"fe9d5501199de618", X"edcf14b4d7ba8180"),
        (X"827af902cd859b23", X"75bfe2cce6c283f1"),
        (X"d8a8c2aaa0e7b685", X"0b8a71febbd7962f"),
        (X"3edd8d0cc4407d2c", X"f8ca4d7a4b4b9e8a"),
        (X"7fd9c13afec846a2", X"f1be90d1adb8f5f8"),
        (X"1d57f851f1175f6f", X"4017e5e578b2b1da"),
        (X"9be255cc6f3e2fd1", X"cb65a286ff70fe4a"),
        (X"4a880453f3fc658d", X"874656316994f261"),
        (X"fda53b04a3987612", X"fc11b5479d19150f"),
        (X"1cbb4fd27f3bd913", X"71b92e68c8bebd0d"),
        (X"68b4c9b977d41fa0", X"1529977556d16376"),
        (X"0bdc40947b43c0b4", X"76b64e3d2a9f32d7"),
        (X"dbf17b83845b268d", X"bf248aa839385465"),
        (X"9f97ed5916776b06", X"633ca2734565881f"),
        (X"dfb91da38950ebf0", X"efee8dd52aa378f8"),
        (X"63a48906dc1947df", X"54a14a45eace37c4"),
        (X"c95e4742e4814c61", X"1c6f8ab2f3292da5"),
        (X"d93075a62d42b0d6", X"94c35440531e3f4e"),
        (X"1f9e759768e597c0", X"1a45ef493a754398"),
        (X"673a145a53cf94ff", X"4048a269ae92d66e"),
        (X"2c1fcaa0090e2218", X"5bc3558dd9d2722b"),
        (X"720e06fc3ab6cf68", X"80273c525e269746"),
        (X"2a0a70d2ee437855", X"cdeb6273d27f5b4f"),
        (X"fb968ddef9bdbe5d", X"f316f7880f64a1e7"),
        (X"be34002f5231d251", X"9c19dd6254b4e977"),
        (X"22de470fee383c5c", X"be7d9a637f9d7e35"),
        (X"f3cf282952f67e4a", X"a11a0e31a6b48a7a"),
        (X"3e04ba1ca6232edc", X"00c6ab9a7fc14d3e"),
        (X"e3e0f332cdbc7f0e", X"711a86cff98ec788"),
        (X"d9bef4ac231d8011", X"e16e8d5a9ee1d0c6"),
        (X"0a499dfd2ccd6350", X"10c84e4e19166d7f"),
        (X"42db76ef773c38ce", X"4ec62875da1fec41"),
        (X"56557e5247908701", X"1fa687abfbda4d15"),
        (X"a4daf3a7c6972aba", X"8e847d066ae41493"),
        (X"e7681c4b715da00c", X"ab58e1b571cb4391"),
        (X"c2d672510b812011", X"70a0a9af1ca59b9b"),
        (X"9955064a7c598e54", X"3aff46b296b9a7e3"),
        (X"4f3e05500c6209df", X"f6c530e34872be5f"),
        (X"7539bddad3d945e4", X"ca48773df186582d"),
        (X"636287313b9b100e", X"f0036db773c85d9a"),
        (X"891ac8406e42266e", X"2cf2b6d7bfe5b39c"),
        (X"e9b89414097b0014", X"21eaebb1d2cbf83e"),
        (X"9b8c9bcb59801dc1", X"b212d94fc40a2540"),
        (X"50e64abbc9ca7bb3", X"9f97316e8396f333"),
        (X"6604164de712d1d6", X"bcc54502d1d12444"),
        (X"d1288263aca828b0", X"b47d9c9064371b45"),
        (X"6be5ac65cfd82b4d", X"b5f56b02d161e2c5"),
        (X"a64e54730490f2e6", X"ad2138ba1f5f0f42"),
        (X"c391e47b63c7ab89", X"6238df14eeee3c08"),
        (X"3cc27767dde132ab", X"951dbe9e9f336127"),
        (X"b28c5444dfc6d3db", X"bef769855e4951a3"),
        (X"da42a21ccd6e59bc", X"d1ac5e19ee0e8a80"),
        (X"3a0a0fe6f3fccdea", X"0e47a5740848c68b"),
        (X"48b32eb1e7a0b6e8", X"4e4a3a3c2e25541d"),
        (X"b08f925fef29cbfd", X"46cdcae66124d21b"),
        (X"675a59c472839109", X"4d24e4a46e750770"),
        (X"68b969399316d450", X"ae3cdad581cccc98"),
        (X"9b982f7a114f93ff", X"05e73b4ae78c35b5"),
        (X"42d899db25877d61", X"1d27ab8e12e7f50a"),
        (X"7ab2e8e907c3af0a", X"dc9861a4121f7059"),
        (X"c69906e08572fdee", X"03811feab1488375"),
        (X"a53a42e2c641a374", X"12f098b7f74c0799"),
        (X"c891ec0025fa9bcd", X"8e2e893927caab0e"),
        (X"718b1b58f2bc5fe6", X"944c4ee754bfba13"),
        (X"1237c3fbb80983b8", X"bce7c8cc9c9d3cf4"),
        (X"d29e66c6ecff36a1", X"d8b7526b2b038ac3"),
        (X"8151ad6f4fabdab3", X"235e33186ad7df8d"),
        (X"ef481c75456b4b07", X"8d5f755823b09e4a"),
        (X"8c8768869a366c74", X"0f39e0dd8924f5ac"),
        (X"914c9f05da8228cd", X"96a018e8bf981239"),
        (X"f9ab13ad19280f35", X"1a298ffe10615636"),
        (X"e57f610d11879ce9", X"07bd4b46d23b7674"),
        (X"ebee359b46a762b3", X"46317e93851b943b"),
        (X"e905506e294e8253", X"ef16c5699faa8b64"),
        (X"38945da34025924a", X"d760eb5574225f5b"),
        (X"4b8a8cee2911bbbc", X"92237ad9905f642b"),
        (X"bc8aa1e206ff586e", X"b128d4f83f03aa43"),
        (X"61fd28f4a3ae5d78", X"b9ee3c785ae35b94"),
        (X"4d79f28947b773f3", X"92f1ca1318a2626c"),
        (X"153974bb7bbddee3", X"6d216bad9ddd8ff7"),
        (X"e1aa98eb6076d664", X"ed9cc8b4874a7ffa"),
        (X"c06fb82079c3e045", X"7e87bf42d0e76bd6"),
        (X"823483bd0a62c9d3", X"9663e6414d615a82"),
        (X"c06339fd566e2e6b", X"6620a3e39ca5619d"),
        (X"e0f3eb9abe01e0af", X"7280ef81f81a4311"),
        (X"915955a637a46c3e", X"b22fa7abfad22e27"),
        (X"b3afd6a96756bc45", X"e9941792efa9284b"),
        (X"e09011e3958af13b", X"e43fd9289bb4d3e2"),
        (X"b356aab276c7e612", X"c36876c99831f1c3"),
        (X"632a542e849d9075", X"7d6aa319f30c90b4"),
        (X"a0d6ea9cdd80fbd2", X"742eddd672a0b2de"),
        (X"b25a77a19b830151", X"66beeca23bb98b1a"),
        (X"67d4f746deb2a406", X"1f7a8c48d506068e"),
        (X"e50df3e868361bca", X"c051b1d8efe3b2bd"),
        (X"ef836e90a73355a9", X"9ba7ac12f7d241ff"),
        (X"9d2a544840d4c050", X"1bd053e7732b54fd"),
        (X"a273633845ae17d4", X"74cbcf3beb5f791f"),
        (X"3ccb8bd0865d4d16", X"16111d2bca923e60"),
        (X"e15011f34261f7d8", X"f2fd7b85a7e4dd22"),
        (X"c297433100e1ae78", X"7e6c1a067bd843cb"),
        (X"543d2324318ad74b", X"bdd92332456c3ef1"),
        (X"648ea461e0700a7b", X"7077506c3157c9d6"),
        (X"fd3a3578c0ef4905", X"1da3896932c92483"),
        (X"9fce7fa40c44533a", X"973bc33e790a13c6"),
        (X"4caad1709cfcdc15", X"da5b6b7509cbab95"),
        (X"80b93372505a4f56", X"145f0bc7e2d5b118"),
        (X"5e4882c203e18413", X"585025dae90a2c07"),
        (X"1ecfb22bfbe7f700", X"80b5a8c89e73e281"),
        (X"cda38ad10c8624cd", X"a9a3a5d58862ef69"),
        (X"86ca132e9217aac1", X"51732dd5144650ab"),
        (X"c00a833bd85bb049", X"c2543adbdc3d8d9a"),
        (X"38549b24f1bdc1e9", X"ee2711f7283e9008"),
        (X"55071c0fcf5bdc12", X"fb9620e86745be19"),
        (X"8b375b15d319a1a9", X"c49f542348df0f18"),
        (X"1398f3d65e127a92", X"ef2dfec0bea287b7"),
        (X"cc597d61b8da15e4", X"655ed0b2b6058d59"),
        (X"0429e6dbf56cc635", X"7bff40d2015e3d8f"),
        (X"d5a6a1d1e4c275be", X"61e3abdf3847e6ec"),
        (X"681a62911a655a40", X"37492e0a9df34df9"),
        (X"ad1e34d963f834cd", X"1c96eff8259c6c07"),
        (X"3baf3053810b0d5c", X"02094a16c5d741e3"),
        (X"7eb48dc3aa56a8b9", X"84e027a241536eac"),
        (X"b5c2e72a51561448", X"6490f942d8220ccb"),
        (X"495d627a845e50a6", X"4076ba710efc4ef9"),
        (X"5322d8f92edaf8d6", X"e08393213fcb3c3d"),
        (X"bd8476985f8ae9c3", X"f087221eb3464403"),
        (X"733b0613838f2403", X"30ff01ee97a1fd08"),
        (X"71ba525081733c5f", X"0b609841224f980d"),
        (X"ae84b7291b39d351", X"a06bc3ad8585b211"),
        (X"eba069f745c41e91", X"0d43333c7000436f"),
        (X"adf25f80b6b8de4c", X"ec2f18886456f695"),
        (X"7a036dfc09e14c6d", X"75555c9d1e7ccfdd"),
        (X"883b0acde25c7c18", X"4cd9e6d4bdcfc872"),
        (X"4868e8f6d19e2aa5", X"922798d0b87da700"),
        (X"8378161f15a0fa17", X"c77597ffe1232eeb"),
        (X"7f15cd0929b4f37a", X"7a92c76ae0858bea"),
        (X"cdc6a6625b6a6906", X"38d3250733f2135e"),
        (X"a16fd1c0ae7160e1", X"bf04af4a1dd111e8"),
        (X"4b72c11bd7c22293", X"9995859466751ef2"),
        (X"5dbbf033b8aed5a8", X"fd4c19dbd4a6cb80"),
        (X"a2193cf6518eadc3", X"b55a60175e157b54"),
        (X"29dce38dc1901257", X"a20c31592ad6c32c"),
        (X"749ece426dca43a5", X"10f565d7e089174e"),
        (X"88fdf085c68fada7", X"d610ee936833b972"),
        (X"7a097fb72745acb8", X"234056819095d693"),
        (X"d7cbe2a19dfe55cd", X"d43db72b8f9d4dc8"),
        (X"59024bae45f6a064", X"6f4fb2dd730ba455"),
        (X"6689c5efa8b4ed33", X"b298c69a16bf387c"),
        (X"741e078acfcf74a5", X"21347219c9267bb1"),
        (X"8cb984909ea305bb", X"e4b9846d01c7db83"),
        (X"b83994ebbe9a1b42", X"071487aedcf22e95"),
        (X"a72a2b0664499a34", X"da3b5dca7f456b95"),
        (X"73a13b6c25a9b921", X"9a84619ef3c8fc1a"),
        (X"a0b68abfa6538c91", X"d3f834e4c0b7ed78"),
        (X"1c03db123db07b47", X"7a8558d6c2565a4a"),
        (X"7bdd161a50c0a36b", X"cc27f1ca5c02411e"),
        (X"0950335041243fc7", X"4ffa76be2c66148d"),
        (X"87c6b714242e3acd", X"0318a7f2b3e73234"),
        (X"e876b8c0b904ecd9", X"27599699bd4194a5"),
        (X"13752f1e1fd14383", X"66b9f67f7d1553a3"),
        (X"e87b931be1767e56", X"12a098053f42404d"),
        (X"cb8e98b861775a46", X"cee8e3e2a7ee3b2e"),
        (X"a7a421b47814f6f3", X"dbada417f5a8f8c6"),
        (X"59e1a963ceae454a", X"1163dff4601899fc"),
        (X"802f809221137329", X"7a589e9488ca47d1"),
        (X"792192a7f2ba8571", X"27f300a02c3e956e"),
        (X"801c7ada922385fa", X"f044f3d37fd572a8"),
        (X"ffe9ac1e35dde2df", X"9e59c6ef24403740"),
        (X"6e622ae82ce02785", X"7dfb06a058a3a4fc"),
        (X"c2f314c9e0928482", X"4ea4ee1666c6dc9f"),
        (X"faa58877f29b80ba", X"781a807d23a4cffb"),
        (X"2fdd8fa725898d12", X"ba2c9860b48104c2"),
        (X"71d10395d235cb4c", X"8ab642223e004e25"),
        (X"7c53a62918bc860b", X"fa0a7af8239672fd"),
        (X"15afac4b39812f49", X"8fe1e8fded846994"),
        (X"a4bc60c76311a359", X"24d8b59d42034fbe"),
        (X"00a4b5d9f26b4058", X"6a4899f49463f513"),
        (X"83e28516856b839b", X"1ff98bdd88d53589"),
        (X"e718847754d4c1ed", X"988a7afd852bd5a0"),
        (X"4a5f3a91f3a1efe5", X"9d6e535c4873ea00"),
        (X"7bdb0dd68c44f3c1", X"e5da9b7c53d68a14"),
        (X"5f8bcc5a39b79f85", X"1728dc9c81e3714c"),
        (X"1f515523eb87abe3", X"6db77cbf46ed430c"),
        (X"71ab3e5ef18cf970", X"0b4476f234f90ed9"),
        (X"f7ebdd942742d8dd", X"d94cb144e88167cc"),
        (X"65ecdca06f28972e", X"f14cb28ea50fd035"),
        (X"0ad9d0e2460c5107", X"dde87b33571ed90a"),
        (X"0fc4df39da176044", X"9e5d23494064c141"),
        (X"f58af2bec0fc9583", X"65596b68156562ce"),
        (X"3168d4754d826fa4", X"15c1fbbade1a0f5a"),
        (X"0f949a5fbecd8185", X"02816dc90cec1bcf"),
        (X"e3b4e2c6390a0d47", X"6ce71801ef47d3f5"),
        (X"1e55fd6c8b57fb42", X"0502437f54c3867b"),
        (X"e1f38b6267bfb38a", X"8a093bcf5c04e18c"),
        (X"03f65bb9a2b44991", X"13f5cf38ade0b6ad"),
        (X"fa74abc7aa914de5", X"743e64daca567487"),
        (X"d0e2a5fc1389a72a", X"070f03a8613c8b9b"),
        (X"f461e326b9a98239", X"50403218e08d40a4"),
        (X"c3061b3b9a419bbc", X"3d66c4727863c242"),
        (X"2d893a9699d255a1", X"5fcaef7895f8a371"),
        (X"2b78a209e5de9dd1", X"728750fdbc3ec91e"),
        (X"37267014bf7978b1", X"8817b70bae866cc5"),
        (X"1f107b009ee4c216", X"c18b60fc75ff0d4c"),
        (X"628d66f42cdda960", X"674edd73e7285dc1"),
        (X"fe1318d97c75fc5c", X"3e54989ebb05a2db"),
        (X"d16897f0068a9012", X"455ce4c883aebd21"),
        (X"43eb2c3af7cf053b", X"d3f3311d54d5ea64"),
        (X"44155f5b6de2f6ae", X"0b0d1517663bb0e7"),
        (X"a78efcc86a9c4a16", X"7e362c54931a7f94"),
        (X"8877bbd4075c44bc", X"abde482e59056093"),
        (X"53b095ebf1079a0c", X"7533425719f712b0"),
        (X"47778c482332817a", X"9f289f061ca48fef"),
        (X"a770ab1a665b06c9", X"c13efa4fe60f6d46"),
        (X"db8d0b95c2ccc208", X"4b3da2240c030bab"),
        (X"7852800f89d16c16", X"18352c69f8198de5"),
        (X"9e7b87581d9ed913", X"8e0bb64f51314914"),
        (X"3b78d7321d7a43fb", X"1e1167d9715eaa70"),
        (X"4f92fc82ced2937c", X"9a728b7d9df31383"),
        (X"6fc8b7d7343b1cd4", X"420a33145969b3f7"),
        (X"873acf362488c650", X"be736d037e4909c3"),
        (X"f09640918320a6ba", X"eee1dea4549a84ed"),
        (X"17bb4df412d67f1d", X"e10b57443a616159"),
        (X"8e9534d8dd84356c", X"1c9b4460d589b6c7"),
        (X"eb410933c76c3e88", X"2ea72747365c54e8"));
end package;

