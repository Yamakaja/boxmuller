library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package pp_fcn_rom_pkg is

    type log_coeff_table_t is array(0 to 255) of std_logic_vector(67 downto 0);
    constant LOG_COEFF_TABLE_DATA : log_coeff_table_t := (
        "10000000100000011111111111111111100110000000000000000000000000000001",
        "10000001100000011111111000000001100110000000001111111110000000010110",
        "10000010011110011111110000000111100010000000011111111000000010101010",
        "10000011011100011111101000010001011010000000101111101110001000111100",
        "10000100011001011111100000011111001000000000111111100000010101000110",
        "10000101010101011111011000110000101010000001001111001110101001000101",
        "10000110010001011111010001000101111110000001011110111001000110110001",
        "10000111001100011111001001011111000000000001101110011111110000000011",
        "10001000000111011111000001111011110000000001111110000010100110110001",
        "10001001000000011110111010011100001000000010001101100001101100110010",
        "10001001111001011110110011000000001000000010011100111101000011111000",
        "10001010110010011110101011100111101010000010101100010100101101110110",
        "10001011101001011110100100010010110000000010111011101000101100011111",
        "10001100100001011110011101000001010100000011001010111001000001100010",
        "10001101010111011110010101110011010100000011011010000101101110101111",
        "10001110001101011110001110101000110000000011101001001110110101110010",
        "10001111000011011110000111100001100010000011111000010100011000011000",
        "10001111110111011110000000011101101010000100000111010110011000001110",
        "10010000101011011101111001011101000110000100010110010100110110111100",
        "10010001011111011101110010011111110010000100100101001111110110001100",
        "10010010010010011101101011100101101100000100110100000111010111100110",
        "10010011000101011101100100101110110100000101000010111011011100110000",
        "10010011110111011101011101111011000100000101010001101100000111010000",
        "10010100101000011101010111001010011110000101100000011001011000101011",
        "10010101011001011101010000011100111100000101101111000011010010100011",
        "10010110001001011101001001110010011110000101111101101001110110011100",
        "10010110111001011101000011001011000010000110001100001101000101110110",
        "10010111101001011100111100100110100110000110011010101101000010010010",
        "10011000011000011100110110000101000110000110101001001001101101001111",
        "10011001000110011100101111100110100010000110110111100011001000001011",
        "10011001110100011100101001001010111000000111000101111001010100100100",
        "10011010100001011100100010110010000110000111010100001100010011110110",
        "10011011001110011100011100011100001010000111100010011100000111011100",
        "10011011111011011100010110001001000000000111110000101000110000110000",
        "10011100100111011100001111111000101010000111111110110010010001001101",
        "10011101010010011100001001101011000010001000001100111000101010001010",
        "10011101111101011100000011100000001010001000011010111011111100111111",
        "10011110101000011011111101010111111110001000101000111100001011000010",
        "10011111010010011011110111010010011100001000110110111001010101101011",
        "10011111111100011011110001001111100100001001000100110011011110001101",
        "10100000100110011011101011001111010010001001010010101010100101111100",
        "10100001001111011011100101010001101000001001100000011110101110001101",
        "10100001110111011011011111010110100000001001101110001111111000010000",
        "10100010011111011011011001011101111010001001111011111110000101011001",
        "10100011000111011011010011100111110110001010001001101001010110110111",
        "10100011101110011011001101110100010000001010010111010001101101111010",
        "10100100010101011011001000000011001000001010100100110111001011110010",
        "10100100111100011011000010010100011100001010110010011001110001101101",
        "10100101100010011010111100101000001010001010111111111001100000111000",
        "10100110001000011010110110111110010010001011001101010110011010100001",
        "10100110101110011010110001010110110000001011011010110000011111110100",
        "10100111010011011010101011110001100100001011101000000111110001111011",
        "10100111110111011010100110001110101110001011110101011100010010000001",
        "10101000011100011010100000101110001010001100000010101110000001010001",
        "10101001000000011010011011001111111000001100001111111101000000110011",
        "10101001100100011010010101110011110100001100011101001001010001101111",
        "10101010000111011010010000011010000010001100101010010010110101001111",
        "10101010101010011010001011000010011100001100110111011001101100010111",
        "10101011001101011010000101101101000010001101000100011101111000010000",
        "10101011101111011010000000011001110010001101010001011111011001111110",
        "10101100010001011001111011001000101100001101011110011110010010100111",
        "10101100110011011001110101111001101110001101101011011010100011001111",
        "10101101010100011001110000101100110110001101111000010100001100111010",
        "10101101110101011001101011100010000110001110000101001011010000101011",
        "10101110010110011001100110011001011000001110010001111111101111100100",
        "10101110110110011001100001010010101110001110011110110001101010100111",
        "10101111010111011001011100001110000110001110101011100001000010110110",
        "10101111110110011001010111001011011110001110111000001101111001010000",
        "10110000010110011001010010001010110110001111000100111000001110110111",
        "10110000110101011001001101001100001100001111010001100000000100101001",
        "10110001010100011001001000001111100000001111011110000101011011100110",
        "10110001110011011001000011010100110000001111101010101000010100101011",
        "10110010010001011000111110011011111010001111110111001000110000110111",
        "10110010110000011000111001100100111100010000000011100110110001000110",
        "10110011001101011000110100101111111010010000010000000010010110010101",
        "10110011101011011000101111111100101110010000011100011011100001100000",
        "10110100001000011000101011001011011000010000101000110010010011100010",
        "10110100100101011000100110011011111000010000110101000110101101011000",
        "10110101000010011000100001101110001100010001000001011000101111111010",
        "10110101011111011000011101000010010010010001001101101000011100000011",
        "10110101111011011000011000011000001100010001011001110101110010101100",
        "10110110010111011000010011101111110110010001100110000000110100101110",
        "10110110110011011000001111001001010010010001110010001001100011000001",
        "10110111001111011000001010100100011100010001111110001111111110011110",
        "10110111101010011000000110000001010100010010001010010100000111111100",
        "10111000000101011000000001011111111010010010010110010110000000010001",
        "10111000100000010111111101000000001100010010100010010101101000010100",
        "10111000111010010111111000100010001010010010101110010011000000111011",
        "10111001010101010111110100000101110010010010111010001110001010111011",
        "10111001101111010111101111101011000010010011000110000111000111001001",
        "10111010001001010111101011010001111100010011010001111101110110011011",
        "10111010100011010111100110111010011110010011011101110010011001100011",
        "10111010111100010111100010100100100110010011101001100100110001010101",
        "10111011010101010111011110010000010110010011110101010100111110100110",
        "10111011101110010111011001111101101000010100000001000011000010000110",
        "10111100000111010111010101101100100000010100001100101110111100101010",
        "10111100100000010111010001011100111100010100011000011000101111000010",
        "10111100111000010111001101001110111000010100100100000000011010000000",
        "10111101010000010111001001000010011000010100101111100101111110010101",
        "10111101101000010111000100110111011000010100111011001001011100110010",
        "10111110000000010111000000101101110110010101000110101010110110000111",
        "10111110011000010110111100100101110110010101010010001010001011000100",
        "10111110101111010110111000011111010100010101011101100111011100010111",
        "10111111000110010110110100011010001110010101101001000010101010110001",
        "10111111011101010110110000010110100110010101110100011011110110111111",
        "10111111110100010110101100010100011010010101111111110011000001110001",
        "11000000001011010110101000010011101010010110001011001000001011110011",
        "11000000100001010110100100010100010010010110010110011011010101110011",
        "11000000111000010110100000010110010110010110100001101100100000011110",
        "11000001001110010110011100011001110100010110101100111011101100100010",
        "11000001100100010110011000011110101000010110111000001000111010101010",
        "11000001111001010110010100100100110100010111000011010100001011100010",
        "11000010001111010110010000101100011000010111001110011101011111110111",
        "11000010100100010110001100110101010010010111011001100100111000010010",
        "11000010111001010110001000111111100000010111100100101010010101100000",
        "11000011001110010110000101001011000100010111101111101101111000001010",
        "11000011100011010110000001010111111100010111111010101111100000111011",
        "11000011111000010101111101100110001000011000000101101111010000011101",
        "11000100001101010101111001110101100110011000010000101101000111011010",
        "11000100100001010101110110000110010110011000011011101001000110011010",
        "11000100110101010101110010011000011000011000100110100011001110000111",
        "11000101001001010101101110101011101010011000110001011011011111001000",
        "11000101011101010101101011000000001100011000111100010001111010000111",
        "11000101110001010101100111010101111110011001000111000110011111101011",
        "11000110000100010101100011101101000000011001010001111001010000011100",
        "11000110011000010101100000000101010000011001011100101010001101000001",
        "11000110101011010101011100011110101100011001100111011001010110000001",
        "11000110111110010101011000111001010110011001110010000110101100000011",
        "11000111010001010101010101010101001100011001111100110010001111101101",
        "11000111100100010101010001110010010000011010000111011100000001100101",
        "11000111110111010101001110010000011100011010010010000100000010010001",
        "11001000001001010101001010101111110100011010011100101010010010010110",
        "11001000011011010101000111010000011000011010100111001110110010011010",
        "11001000101110010101000011110010000100011010110001110001100011000010",
        "11001001000000010101000000010100111000011010111100010010100100110010",
        "11001001010010010100111100111000110110011011000110110001111000001111",
        "11001001100100010100111001011101111010011011010001001111011101111100",
        "11001001110101010100110110000100000110011011011011101011010110011101",
        "11001010000111010100110010101011011010011011100110000101100010010110",
        "11001010011000010100101111010011110100011011110000011110000010001011",
        "11001010101010010100101011111101010010011011111010110100110110011101",
        "11001010111011010100101000100111110110011100000101001001111111110001",
        "11001011001100010100100101010011100000011100001111011101011110101000",
        "11001011011101010100100010000000001100011100011001101111010011100100",
        "11001011101101010100011110101101111110011100100011111111011111000111",
        "11001011111110010100011011011100110010011100101110001110000001110100",
        "11001100001111010100011000001100101000011100111000011010111100001011",
        "11001100011111010100010100111101100000011101000010100110001110101110",
        "11001100101111010100010001101111011010011101001100101111111001111110",
        "11001100111111010100001110100010010110011101010110110111111110011011",
        "11001101010000010100001011010110010010011101100000111110011100100101",
        "11001101011111010100001000001011001110011101101011000011010100111110",
        "11001101101111010100000101000001001010011101110101000110101000000101",
        "11001101111111010100000001111000000100011101111111001000010110011001",
        "11001110001111010011111110101111111110011110001001001000100000011010",
        "11001110011110010011111011101000110110011110010011000111000110101000",
        "11001110101101010011111000100010101100011110011101000100001001100010",
        "11001110111101010011110101011101100000011110100110111111101001100101",
        "11001111001100010011110010011001010000011110110000111001100111010010",
        "11001111011011010011101111010101111100011110111010110010000011000110",
        "11001111101010010011101100010011100110011111000100101000111101011111",
        "11001111111000010011101001010010001010011111001110011110010110111100",
        "11010000000111010011100110010001101010011111011000010010001111111010",
        "11010000010110010011100011010010000100011111100010000100101000110111",
        "11010000100100010011100000010011011010011111101011110101100010001111",
        "11010000110011010011011101010101101000011111110101100100111100100001",
        "11010001000001010011011010011000110010011111111111010010111000001000",
        "11010001001111010011010111011100110010100000001000111111010101100010",
        "11010001011101010011010100100001101110100000010010101010010101001011",
        "11010001101011010011010001100111100000100000011100010011110111011111",
        "11010001111001010011001110101110001010100000100101111011111100111011",
        "11010010000111010011001011110101101110100000101111100010100101111010",
        "11010010010101010011001000111110000110100000111001000111110010111000",
        "11010010100010010011000110000111010110100001000010101011100100010000",
        "11010010110000010011000011010001011110100001001100001101111010011110",
        "11010010111101010011000000011100011010100001010101101110110101111101",
        "11010011001010010010111101101000001100100001011111001110010111001000",
        "11010011011000010010111010110100110100100001101000101100011110011001",
        "11010011100101010010111000000010010000100001110010001001001100001011",
        "11010011110010010010110101010000100010100001111011100100100000111001",
        "11010011111111010010110010011111101000100010000100111110011100111100",
        "11010100001100010010101111101111100000100010001110010111000000101111",
        "11010100011000010010101101000000001100100010010111101110001100101011",
        "11010100100101010010101010010001101100100010100001000100000001001010",
        "11010100110010010010100111100011111110100010101010011000011110100110",
        "11010100111110010010100100110111000100100010110011101011100101010111",
        "11010101001011010010100010001010111010100010111100111101010101110111",
        "11010101010111010010011111011111100010100011000110001101110000100000",
        "11010101100011010010011100110100111100100011001111011100110101101001",
        "11010101101111010010011010001011001000100011011000101010100101101011",
        "11010101111100010010010111100010000100100011100001110111000000111111",
        "11010110001000010010010100111001110000100011101011000010000111111101",
        "11010110010100010010010010010010001100100011110100001011111010111101",
        "11010110011111010010001111101011011000100011111101010100011010010111",
        "11010110101011010010001101000101010100100100000110011011100110100011",
        "11010110110111010010001010011111111110100100001111100001011111111000",
        "11010111000010010010000111111011011000100100011000100110000110101111",
        "11010111001110010010000101010111100000100100100001101001011011011110",
        "11010111011010010010000010110100010110100100101010101011011110011101",
        "11010111100101010010000000010001111010100100110011101100010000000010",
        "11010111110000010001111101110000001100100100111100101011110000100101",
        "11010111111011010001111011001111001100100101000101101010000000011100",
        "11011000000111010001111000101110111000100101001110100110111111111101",
        "11011000010010010001110110001111010000100101010111100010101111100000",
        "11011000011101010001110011110000010110100101100000011101001111011010",
        "11011000101000010001110001010010000110100101101001010110100000000010",
        "11011000110011010001101110110100100100100101110010001110100001101101",
        "11011000111101010001101100010111101100100101111011000101010100110010",
        "11011001001000010001101001111011100000100110000011111010111001100110",
        "11011001010011010001100111100000000000100110001100101111010000011111",
        "11011001011110010001100101000101001000100110010101100010011001110010",
        "11011001101000010001100010101010111100100110011110010100010101110100",
        "11011001110011010001100000010001011100100110100111000101000100111011",
        "11011001111101010001011101111000100100100110101111110100100111011011",
        "11011010000111010001011011100000010110100110111000100010111101101010",
        "11011010010010010001011001001000110000100111000001010000000111111100",
        "11011010011100010001010110110001110100100111001001111100000110100110",
        "11011010100110010001010100011011100010100111010010100110111001111101",
        "11011010110000010001010010000101111000100111011011010000100010010100",
        "11011010111010010001001111110000110110100111100011111001000000000000",
        "11011011000100010001001101011100011100100111101100100000010011010101",
        "11011011001110010001001011001000101010100111110101000110011100100111",
        "11011011011000010001001000110101011110100111111101101011011100001001",
        "11011011100001010001000110100010111100101000000110001111010010010001",
        "11011011101011010001000100010001000000101000001110110001111111010000",
        "11011011110101010001000001111111101010101000010111010011100011011011",
        "11011011111110010000111111101110111100101000011111110011111111000110",
        "11011100001000010000111101011110110100101000101000010011010010100010",
        "11011100010001010000111011001111010000101000110000110001011110000100",
        "11011100011011010000111001000000010100101000111001001110100001111110",
        "11011100100100010000110110110001111110101001000001101010011110100011",
        "11011100101101010000110100100100001100101001001010000101010100000111",
        "11011100110111010000110010010111000000101001010010011111000010111011",
        "11011101000000010000110000001010011010101001011010110111101011010010",
        "11011101001001010000101101111110011000101001100011001111001101011111",
        "11011101010010010000101011110010111010101001101011100101101001110100",
        "11011101011011010000101001101000000000101001110011111011000000100011",
        "11011101100100010000100111011101101010101001111100001111010001111110",
        "11011101101101010000100101010011111000101010000100100010011110011000",
        "11011101110110010000100011001010101010101010001100110100100110000001",
        "11011101111111010000100001000010000000101010010101000101101001001100",
        "11011110000111010000011110111001111000101010011101010101101000001011",
        "11011110010000010000011100110010010100101010100101100100100011001111",
        "11011110011001010000011010101011010010101010101101110010011010101001",
        "11011110100001010000011000100100110010101010110101111111001110101011",
        "11011110101010010000010110011110110110101010111110001010111111100110",
        "11011110110010010000010100011001011100101011000110010101101101101011",
        "11011110111011010000010010010100100010101011001110011111011001001100",
        "11011111000011010000010000010000001100101011010110101000000010011000",
        "11011111001011010000001110001100010110101011011110101111101001100001",
        "11011111010100010000001100001001000010101011100110110110001110111000",
        "11011111011100010000001010000110010000101011101110111011110010101110",
        "11011111100100010000001000000011111110101011110111000000010101010010",
        "11011111101100010000000110000010001100101011111111000011110110110101",
        "11011111110100010000000100000000111100101100000111000110010111101000",
        "11011111111100010000000010000000001100101100001111000111110111111011"
    );
    
    type sqrt_coeff_table_t is array(0 to 127) of std_logic_vector(31 downto 0);
    constant SQRT_COEFF_TABLE_DATA : sqrt_coeff_table_t := (
        "00111111110000000000000000000001",
        "00111111010000000000011111111001",
        "00111110110010000000111111100001",
        "00111110010100000001011110111010",
        "00111101110110000001111110000101",
        "00111101011010000010011101000000",
        "00111100111110000010111011101101",
        "00111100100010000011011010001101",
        "00111100001000000011111000011110",
        "00111011101110000100010110100010",
        "00111011010100000100110100011010",
        "00111010111010000101010010000100",
        "00111010100010000101101111100001",
        "00111010001010000110001100110011",
        "00111001110010000110101001111000",
        "00111001011010000111000110110001",
        "00111001000100000111100011011110",
        "00111000101100001000000000000000",
        "00111000010110001000011100010111",
        "00111000000000001000111000100011",
        "00110111101100001001010100100100",
        "00110111010110001001110000011010",
        "00110111000010001010001100000110",
        "00110110101110001010100111101000",
        "00110110011010001011000010111111",
        "00110110000110001011011110001101",
        "00110101110100001011111001010001",
        "00110101100000001100010100001011",
        "00110101001110001100101110111100",
        "00110100111100001101001001100011",
        "00110100101010001101100100000010",
        "00110100011000001101111110010111",
        "00110100000110001110011000100100",
        "00110011110110001110110010101000",
        "00110011100100001111001100100011",
        "00110011010100001111100110010110",
        "00110011000100010000000000000000",
        "00110010110100010000011001100010",
        "00110010100100010000110010111101",
        "00110010010100010001001100001111",
        "00110010000100010001100101011001",
        "00110001110110010001111110011100",
        "00110001100110010010010111010111",
        "00110001011000010010110000001011",
        "00110001001000010011001000110111",
        "00110000111010010011100001011100",
        "00110000101100010011111001111010",
        "00110000011110010100010010010000",
        "00110000010000010100101010100000",
        "00110000000010010101000010101001",
        "00101111110110010101011010101011",
        "00101111101000010101110010100110",
        "00101111011010010110001010011010",
        "00101111001110010110100010001000",
        "00101111000010010110111001110000",
        "00101110110100010111010001010001",
        "00101110101000010111101000101011",
        "00101110011100011000000000000000",
        "00101110010000011000010111001110",
        "00101110000100011000101110010111",
        "00101101111000011001000101011001",
        "00101101101100011001011100010101",
        "00101101100000011001110011001100",
        "00101101010100011010001001111101",
        "01011010001010011010100000101001",
        "01011001011100011011001101101110",
        "01011000110010011011111010011101",
        "01011000001000011100100110110110",
        "01010111011110011101010010111010",
        "01010110110110011101111110101010",
        "01010110001110011110101010000101",
        "01010101101000011111010101001101",
        "01010101000010100000000000000001",
        "01010100011100100000101010100010",
        "01010011111000100001010100110001",
        "01010011010100100001111110101101",
        "01010010110010100010101000011000",
        "01010010001110100011010001110001",
        "01010001101110100011111010111001",
        "01010001001100100100100011110000",
        "01010000101100100101001100010111",
        "01010000001100100101110100101101",
        "01001111101100100110011100110100",
        "01001111001110100111000100101011",
        "01001110110000100111101100010011",
        "01001110010010101000010011101011",
        "01001101110110101000111010110101",
        "01001101011010101001100001110000",
        "01001100111100101010001000011101",
        "01001100100010101010101110111100",
        "01001100000110101011010101001101",
        "01001011101100101011111011010001",
        "01001011010010101100100001000111",
        "01001010111000101101000110110001",
        "01001010011110101101101100001101",
        "01001010000110101110010001011100",
        "01001001101100101110110110011111",
        "01001001010100101111011011010110",
        "01001000111100110000000000000000",
        "01001000100100110000100100011111",
        "01001000001110110001001000110010",
        "01000111110110110001101100111001",
        "01000111100000110010010000110101",
        "01000111001010110010110100100110",
        "01000110110100110011011000001011",
        "01000110011110110011111011100110",
        "01000110001010110100011110110110",
        "01000101110100110101000001111011",
        "01000101100000110101100100110110",
        "01000101001100110110000111100110",
        "01000100111000110110101010001100",
        "01000100100100110111001100101001",
        "01000100010000110111101110111011",
        "01000011111100111000010001000011",
        "01000011101010111000110011000010",
        "01000011010110111001010100111000",
        "01000011000100111001110110100100",
        "01000010110010111010011000000110",
        "01000010100000111010111001100000",
        "01000010001110111011011010110000",
        "01000001111100111011111011111000",
        "01000001101100111100011100110111",
        "01000001011010111100111101101101",
        "01000001001000111101011110011010",
        "01000000111000111101111110111111",
        "01000000101000111110011111011100",
        "01000000011000111110111111110000",
        "01000000001000111111011111111100"
    );
    
    type trig_coeff_table_t is array(0 to 127) of std_logic_vector(61 downto 0);
    constant TRIG_COEFF_TABLE_DATA : trig_coeff_table_t := (
        "01100100100000000000000000000001111111101110100000000000000001",
        "01100100100000000000110010010001111111000110011111111111110111",
        "01100100011100000001100100100001111110011110011111111111011010",
        "01100100011100000010010110110001111101110110011111111110101000",
        "01100100011000000011001000111111111101010000011111111101100011",
        "01100100010000000011111011001011111100101000011111111100001010",
        "01100100001100000100101101010101111100000000011111111010011110",
        "01100100000100000101011111011011111011011010011111111000011110",
        "01100011111100000110010001011111111010110010011111110110001010",
        "01100011110100000111000011011111111010001010011111110011100011",
        "01100011101100000111110101011001111001100100011111110000100111",
        "01100011100000001000100111001111111000111100011111101101011001",
        "01100011010100001001011001000001111000010110011111101001110110",
        "01100011001000001010001010101101110111101110011111100110000001",
        "01100010111100001010111100010001110111001000011111100001110111",
        "01100010101100001011101101101111110110100000011111011101011011",
        "01100010011100001100011111000111110101111010011111011000101011",
        "01100010001100001101010000010101110101010100011111010011100111",
        "01100001111100001110000001011101110100101100011111001110010000",
        "01100001101000001110110010011011110100000110011111001000100110",
        "01100001010100001111100011010001110011100000011111000010101001",
        "01100001000000010000010011111101110010111010011110111100011001",
        "01100000101100010001000100011111110010010100011110110101110101",
        "01100000011000010001110100110101110001101110011110101110111111",
        "01100000000000010010100101000001110001001000011110100111110101",
        "01011111101000010011010101000011110000100010011110100000011001",
        "01011111010000010100000100110111101111111110011110011000101010",
        "01011110110100010100110100011111101111011000011110010000101000",
        "01011110011100010101100011111011101110110010011110001000010011",
        "01011110000000010110010011001001101110001110011101111111101100",
        "01011101100100010111000010001001101101101000011101110110110010",
        "01011101000100010111110000111011101101000100011101101101100110",
        "01011100101000011000011111011111101100100000011101100100001000",
        "01011100001000011001001101110011101011111100011101011010010111",
        "01011011101000011001111011111001101011011000011101010000010100",
        "01011011001000011010101001101101101010110100011101000101111111",
        "01011010100100011011010111010011101010010000011100111011011001",
        "01011010000100011100000100100111101001101100011100110000100000",
        "01011001100000011100110001101001101001001010011100100101010110",
        "01011000111100011101011110011001101000100110011100011001111010",
        "01011000010100011110001010110111101000000100011100001110001100",
        "01010111110000011110110111000011100111100000011100000010001101",
        "01010111001000011111100010111011100110111110011011110101111101",
        "01010110100000100000001110100001100110011100011011101001011100",
        "01010101111000100000111001110011100101111010011011011100101001",
        "01010101010000100001100100101111100101011000011011001111100110",
        "01010100100100100010001111011001100100111000011011000010010010",
        "01010011111000100010111001101011100100010110011010110100101101",
        "01010011001100100011100011101001100011110110011010100110110111",
        "01010010100000100100001101010001100011010100011010011000110001",
        "01010001110100100100110110100011100010110100011010001010011011",
        "01010001000100100101011111011101100010010100011001111011110101",
        "01010000011000100110001000000001100001110100011001101100111111",
        "01001111101000100110110000001101100001010110011001011101111001",
        "01001110110100100111011000000001100000110110011001001110100011",
        "01001110000100100111111111011101100000011000011000111110111110",
        "01001101010100101000100110100001011111111000011000101111001001",
        "01001100100000101001001101001011011111011010011000011111000101",
        "01001011101100101001110011011011011110111100011000001110110010",
        "01001010111000101010011001010011011110100000010111111110010000",
        "01001010000100101010111110101111011110000010010111101101011111",
        "01001001001100101011100011110001011101100110010111011100011111",
        "01001000011000101100001000011001011101001000010111001011010001",
        "01000111100000101100101100100101011100101100010110111001110101",
        "01000110101000101101010000010111011100010000010110101000001011",
        "01000101110000101101110011101011011011110100010110010110010010",
        "01000100110100101110010110100011011011011010010110000100001100",
        "01000011111100101110111000111111011010111110010101110001111000",
        "01000011000000101111011010111111011010100100010101011111010111",
        "01000010001000101111111100100001011010001010010101001100101001",
        "01000001001100110000011101100101011001110000010100111001101101",
        "01000000010000110000111110001011011001010110010100100110100101",
        "00111111010000110001011110010011011000111110010100010011010000",
        "00111110010100110001111101111101011000100110010011111111101110",
        "00111101010100110010011101000111011000001100010011101100000000",
        "00111100011000110010111011110011010111110100010011011000000110",
        "00111011011000110011011001111111010111011110010011000100000000",
        "00111010011000110011110111101011010111000110010010101111101110",
        "00111001011000110100010100110111010110110000010010011011010001",
        "00111000010100110100110001100011010110011010010010000110101000",
        "00110111010100110101001101101111010110000100010001110001110100",
        "00110110010000110101101001011011010101101110010001011100110101",
        "00110101010000110110000100100101010101011000010001000111101100",
        "00110100001100110110011111001101010101000100010000110010010111",
        "00110011001000110110111001010011010100110000010000011100111001",
        "00110010000100110111010010111001010100011100010000000111010000",
        "00110001000000110111101011111011010100001000001111110001011101",
        "00101111111000111000000100011011010011110110001111011011100001",
        "00101110110100111000011100011001010011100010001111000101011011",
        "00101101101100111000110011110101010011010000001110101111001100",
        "00101100101000111001001010101101010010111110001110011000110100",
        "00101011100000111001100001000001010010101110001110000010010011",
        "00101010011000111001110110110011010010011100001101101011101001",
        "00101001010000111010001011111111010010001100001101010100110110",
        "00101000001000111010100000101001010001111100001100111101111100",
        "00100111000000111010110100101111010001101100001100100110111001",
        "00100101111000111011001000010001010001011110001100001111101111",
        "00100100110000111011011011001101010001001110001011111000011101",
        "00100011100100111011101101100101010001000000001011100001000100",
        "00100010011100111011111111011001010000110010001011001001100100",
        "00100001010000111100010000100111010000100110001010110001111101",
        "00100000000100111100100001010001010000011000001010011010001111",
        "00011110111100111100110001010101010000001100001010000010011011",
        "00011101110000111101000000110011010000000000001001101010100001",
        "00011100100100111101001111101011001111110100001001010010100000",
        "00011011011000111101011101111111001111101010001000111010011010",
        "00011010001100111101101011101011001111100000001000100010001111",
        "00011001000000111101111000110011001111010110001000001001111110",
        "00010111110100111110000101010011001111001100000111110001101000",
        "00010110101000111110010001001101001111000010000111011001001101",
        "00010101011000111110011100100001001110111010000111000000101110",
        "00010100001100111110100111001111001110110010000110101000001010",
        "00010011000000111110110001010111001110101010000110001111100011",
        "00010001110000111110111010110111001110100010000101110110110111",
        "00010000100100111111000011101111001110011100000101011110001000",
        "00001111010100111111001100000011001110010110000101000101010110",
        "00001110001000111111010011101101001110010000000100101100100000",
        "00001100111000111111011010110011001110001010000100010011100111",
        "00001011101100111111100001001111001110000110000011111010101100",
        "00001010011100111111100111000111001110000010000011100001101111",
        "00001001001100111111101100010101001101111110000011001000101111",
        "00001000000000111111110000111101001101111010000010101111101101",
        "00000110110000111111110100111101001101111000000010010110101010",
        "00000101100000111111111000010101001101110100000001111101100101",
        "00000100010100111111111011000111001101110010000001100100011111",
        "00000011000100111111111101010001001101110010000001001011011000",
        "00000001110100111111111110110101001101110000000000110010010000",
        "00000000100100111111111111101111001101110000000000011001001000"
    );

end package;